library verilog;
use verilog.vl_types.all;
entity somador1_vlg_vec_tst is
end somador1_vlg_vec_tst;
